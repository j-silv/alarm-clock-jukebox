-- qsys_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity qsys_system is
	port (
		buttons_external_connection_export    : in  std_logic_vector(1 downto 0) := (others => '0'); --    buttons_external_connection.export
		clk_clk                               : in  std_logic                    := '0';             --                            clk.clk
		hour0_external_connection_export      : out std_logic_vector(7 downto 0);                    --      hour0_external_connection.export
		hour1_external_connection_export      : out std_logic_vector(7 downto 0);                    --      hour1_external_connection.export
		led_alarm_external_connection_export  : out std_logic;                                       --  led_alarm_external_connection.export
		led_piano_external_connection_export  : out std_logic_vector(6 downto 0);                    --  led_piano_external_connection.export
		led_status_external_connection_export : out std_logic_vector(1 downto 0);                    -- led_status_external_connection.export
		minute0_external_connection_export    : out std_logic_vector(7 downto 0);                    --    minute0_external_connection.export
		minute1_external_connection_export    : out std_logic_vector(7 downto 0);                    --    minute1_external_connection.export
		pwm_external_connection_export        : out std_logic;                                       --        pwm_external_connection.export
		reset_reset_n                         : in  std_logic                    := '0';             --                          reset.reset_n
		second0_external_connection_export    : out std_logic_vector(7 downto 0);                    --    second0_external_connection.export
		second1_external_connection_export    : out std_logic_vector(7 downto 0);                    --    second1_external_connection.export
		switches_external_connection_export   : in  std_logic_vector(9 downto 0) := (others => '0')  --   switches_external_connection.export
	);
end entity qsys_system;

architecture rtl of qsys_system is
	component qsys_system_NiosII_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component qsys_system_NiosII_CPU;

	component qsys_system_buttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component qsys_system_buttons;

	component qsys_system_hour0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component qsys_system_hour0;

	component qsys_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component qsys_system_jtag_uart_0;

	component qsys_system_led_alarm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component qsys_system_led_alarm;

	component qsys_system_led_piano is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component qsys_system_led_piano;

	component qsys_system_led_status is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component qsys_system_led_status;

	component qsys_system_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component qsys_system_onchip_memory;

	component pwm_avalon_interface is
		generic (
			clock_divide_reg_init : std_logic_vector(33 downto 0) := "0000000000000000000000000000000000";
			duty_cycle_reg_init   : std_logic_vector(33 downto 0) := "0000000000000000000000000000000000"
		);
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			pwm_out            : out std_logic;                                        -- export
			resetn             : in  std_logic                     := 'X';             -- reset_n
			avalon_chip_select : in  std_logic                     := 'X';             -- chipselect
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write              : in  std_logic                     := 'X';             -- write
			write_data         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read               : in  std_logic                     := 'X';             -- read
			read_data          : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component pwm_avalon_interface;

	component qsys_system_switches is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component qsys_system_switches;

	component qsys_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component qsys_system_sysid_qsys_0;

	component qsys_system_timer_pwm is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component qsys_system_timer_pwm;

	component qsys_system_timer_second is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component qsys_system_timer_second;

	component qsys_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                 : in  std_logic                     := 'X';             -- clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			NiosII_CPU_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			NiosII_CPU_data_master_address                : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			NiosII_CPU_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			NiosII_CPU_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NiosII_CPU_data_master_read                   : in  std_logic                     := 'X';             -- read
			NiosII_CPU_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			NiosII_CPU_data_master_write                  : in  std_logic                     := 'X';             -- write
			NiosII_CPU_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NiosII_CPU_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			NiosII_CPU_instruction_master_address         : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			NiosII_CPU_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			NiosII_CPU_instruction_master_read            : in  std_logic                     := 'X';             -- read
			NiosII_CPU_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			NiosII_CPU_instruction_master_readdatavalid   : out std_logic;                                        -- readdatavalid
			buttons_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			buttons_s1_write                              : out std_logic;                                        -- write
			buttons_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			buttons_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			buttons_s1_chipselect                         : out std_logic;                                        -- chipselect
			hour0_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			hour0_s1_write                                : out std_logic;                                        -- write
			hour0_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hour0_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			hour0_s1_chipselect                           : out std_logic;                                        -- chipselect
			hour1_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			hour1_s1_write                                : out std_logic;                                        -- write
			hour1_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hour1_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			hour1_s1_chipselect                           : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write           : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read            : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect      : out std_logic;                                        -- chipselect
			led_alarm_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			led_alarm_s1_write                            : out std_logic;                                        -- write
			led_alarm_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_alarm_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			led_alarm_s1_chipselect                       : out std_logic;                                        -- chipselect
			led_piano_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			led_piano_s1_write                            : out std_logic;                                        -- write
			led_piano_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_piano_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			led_piano_s1_chipselect                       : out std_logic;                                        -- chipselect
			led_status_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			led_status_s1_write                           : out std_logic;                                        -- write
			led_status_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_status_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			led_status_s1_chipselect                      : out std_logic;                                        -- chipselect
			minute0_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			minute0_s1_write                              : out std_logic;                                        -- write
			minute0_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			minute0_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			minute0_s1_chipselect                         : out std_logic;                                        -- chipselect
			minute1_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			minute1_s1_write                              : out std_logic;                                        -- write
			minute1_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			minute1_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			minute1_s1_chipselect                         : out std_logic;                                        -- chipselect
			NiosII_CPU_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			NiosII_CPU_debug_mem_slave_write              : out std_logic;                                        -- write
			NiosII_CPU_debug_mem_slave_read               : out std_logic;                                        -- read
			NiosII_CPU_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NiosII_CPU_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			NiosII_CPU_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			NiosII_CPU_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			NiosII_CPU_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			onchip_memory_s1_address                      : out std_logic_vector(15 downto 0);                    -- address
			onchip_memory_s1_write                        : out std_logic;                                        -- write
			onchip_memory_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_s1_byteenable                   : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_memory_s1_clken                        : out std_logic;                                        -- clken
			pwm_control_slave_address                     : out std_logic_vector(1 downto 0);                     -- address
			pwm_control_slave_write                       : out std_logic;                                        -- write
			pwm_control_slave_read                        : out std_logic;                                        -- read
			pwm_control_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pwm_control_slave_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			pwm_control_slave_chipselect                  : out std_logic;                                        -- chipselect
			second0_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			second0_s1_write                              : out std_logic;                                        -- write
			second0_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			second0_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			second0_s1_chipselect                         : out std_logic;                                        -- chipselect
			second1_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			second1_s1_write                              : out std_logic;                                        -- write
			second1_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			second1_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			second1_s1_chipselect                         : out std_logic;                                        -- chipselect
			switches_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_write                             : out std_logic;                                        -- write
			switches_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			switches_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			switches_s1_chipselect                        : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address            : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_pwm_s1_address                          : out std_logic_vector(2 downto 0);                     -- address
			timer_pwm_s1_write                            : out std_logic;                                        -- write
			timer_pwm_s1_readdata                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_pwm_s1_writedata                        : out std_logic_vector(15 downto 0);                    -- writedata
			timer_pwm_s1_chipselect                       : out std_logic;                                        -- chipselect
			timer_second_s1_address                       : out std_logic_vector(2 downto 0);                     -- address
			timer_second_s1_write                         : out std_logic;                                        -- write
			timer_second_s1_readdata                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_second_s1_writedata                     : out std_logic_vector(15 downto 0);                    -- writedata
			timer_second_s1_chipselect                    : out std_logic                                         -- chipselect
		);
	end component qsys_system_mm_interconnect_0;

	component qsys_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component qsys_system_irq_mapper;

	component qsys_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component qsys_system_rst_controller;

	component qsys_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component qsys_system_rst_controller_001;

	signal niosii_cpu_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:NiosII_CPU_data_master_readdata -> NiosII_CPU:d_readdata
	signal niosii_cpu_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:NiosII_CPU_data_master_waitrequest -> NiosII_CPU:d_waitrequest
	signal niosii_cpu_data_master_debugaccess                              : std_logic;                     -- NiosII_CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NiosII_CPU_data_master_debugaccess
	signal niosii_cpu_data_master_address                                  : std_logic_vector(19 downto 0); -- NiosII_CPU:d_address -> mm_interconnect_0:NiosII_CPU_data_master_address
	signal niosii_cpu_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- NiosII_CPU:d_byteenable -> mm_interconnect_0:NiosII_CPU_data_master_byteenable
	signal niosii_cpu_data_master_read                                     : std_logic;                     -- NiosII_CPU:d_read -> mm_interconnect_0:NiosII_CPU_data_master_read
	signal niosii_cpu_data_master_write                                    : std_logic;                     -- NiosII_CPU:d_write -> mm_interconnect_0:NiosII_CPU_data_master_write
	signal niosii_cpu_data_master_writedata                                : std_logic_vector(31 downto 0); -- NiosII_CPU:d_writedata -> mm_interconnect_0:NiosII_CPU_data_master_writedata
	signal niosii_cpu_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:NiosII_CPU_instruction_master_readdata -> NiosII_CPU:i_readdata
	signal niosii_cpu_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:NiosII_CPU_instruction_master_waitrequest -> NiosII_CPU:i_waitrequest
	signal niosii_cpu_instruction_master_address                           : std_logic_vector(19 downto 0); -- NiosII_CPU:i_address -> mm_interconnect_0:NiosII_CPU_instruction_master_address
	signal niosii_cpu_instruction_master_read                              : std_logic;                     -- NiosII_CPU:i_read -> mm_interconnect_0:NiosII_CPU_instruction_master_read
	signal niosii_cpu_instruction_master_readdatavalid                     : std_logic;                     -- mm_interconnect_0:NiosII_CPU_instruction_master_readdatavalid -> NiosII_CPU:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_pwm_control_slave_chipselect                  : std_logic;                     -- mm_interconnect_0:pwm_control_slave_chipselect -> pwm:avalon_chip_select
	signal mm_interconnect_0_pwm_control_slave_readdata                    : std_logic_vector(31 downto 0); -- pwm:read_data -> mm_interconnect_0:pwm_control_slave_readdata
	signal mm_interconnect_0_pwm_control_slave_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pwm_control_slave_address -> pwm:address
	signal mm_interconnect_0_pwm_control_slave_read                        : std_logic;                     -- mm_interconnect_0:pwm_control_slave_read -> pwm:read
	signal mm_interconnect_0_pwm_control_slave_write                       : std_logic;                     -- mm_interconnect_0:pwm_control_slave_write -> pwm:write
	signal mm_interconnect_0_pwm_control_slave_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:pwm_control_slave_writedata -> pwm:write_data
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata           : std_logic_vector(31 downto 0); -- NiosII_CPU:debug_mem_slave_readdata -> mm_interconnect_0:NiosII_CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest        : std_logic;                     -- NiosII_CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:NiosII_CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess        : std_logic;                     -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_debugaccess -> NiosII_CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_address -> NiosII_CPU:debug_mem_slave_address
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_read               : std_logic;                     -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_read -> NiosII_CPU:debug_mem_slave_read
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_byteenable -> NiosII_CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_write              : std_logic;                     -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_write -> NiosII_CPU:debug_mem_slave_write
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_writedata -> NiosII_CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	signal mm_interconnect_0_onchip_memory_s1_readdata                     : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_address                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	signal mm_interconnect_0_onchip_memory_s1_byteenable                   : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	signal mm_interconnect_0_onchip_memory_s1_write                        : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	signal mm_interconnect_0_onchip_memory_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	signal mm_interconnect_0_onchip_memory_s1_clken                        : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	signal mm_interconnect_0_switches_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:switches_s1_chipselect -> switches:chipselect
	signal mm_interconnect_0_switches_s1_readdata                          : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal mm_interconnect_0_switches_s1_write                             : std_logic;                     -- mm_interconnect_0:switches_s1_write -> mm_interconnect_0_switches_s1_write:in
	signal mm_interconnect_0_switches_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:switches_s1_writedata -> switches:writedata
	signal mm_interconnect_0_led_piano_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:led_piano_s1_chipselect -> led_piano:chipselect
	signal mm_interconnect_0_led_piano_s1_readdata                         : std_logic_vector(31 downto 0); -- led_piano:readdata -> mm_interconnect_0:led_piano_s1_readdata
	signal mm_interconnect_0_led_piano_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_piano_s1_address -> led_piano:address
	signal mm_interconnect_0_led_piano_s1_write                            : std_logic;                     -- mm_interconnect_0:led_piano_s1_write -> mm_interconnect_0_led_piano_s1_write:in
	signal mm_interconnect_0_led_piano_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_piano_s1_writedata -> led_piano:writedata
	signal mm_interconnect_0_hour0_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:hour0_s1_chipselect -> hour0:chipselect
	signal mm_interconnect_0_hour0_s1_readdata                             : std_logic_vector(31 downto 0); -- hour0:readdata -> mm_interconnect_0:hour0_s1_readdata
	signal mm_interconnect_0_hour0_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hour0_s1_address -> hour0:address
	signal mm_interconnect_0_hour0_s1_write                                : std_logic;                     -- mm_interconnect_0:hour0_s1_write -> mm_interconnect_0_hour0_s1_write:in
	signal mm_interconnect_0_hour0_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:hour0_s1_writedata -> hour0:writedata
	signal mm_interconnect_0_minute0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:minute0_s1_chipselect -> minute0:chipselect
	signal mm_interconnect_0_minute0_s1_readdata                           : std_logic_vector(31 downto 0); -- minute0:readdata -> mm_interconnect_0:minute0_s1_readdata
	signal mm_interconnect_0_minute0_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:minute0_s1_address -> minute0:address
	signal mm_interconnect_0_minute0_s1_write                              : std_logic;                     -- mm_interconnect_0:minute0_s1_write -> mm_interconnect_0_minute0_s1_write:in
	signal mm_interconnect_0_minute0_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:minute0_s1_writedata -> minute0:writedata
	signal mm_interconnect_0_second0_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:second0_s1_chipselect -> second0:chipselect
	signal mm_interconnect_0_second0_s1_readdata                           : std_logic_vector(31 downto 0); -- second0:readdata -> mm_interconnect_0:second0_s1_readdata
	signal mm_interconnect_0_second0_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:second0_s1_address -> second0:address
	signal mm_interconnect_0_second0_s1_write                              : std_logic;                     -- mm_interconnect_0:second0_s1_write -> mm_interconnect_0_second0_s1_write:in
	signal mm_interconnect_0_second0_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:second0_s1_writedata -> second0:writedata
	signal mm_interconnect_0_timer_second_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:timer_second_s1_chipselect -> timer_second:chipselect
	signal mm_interconnect_0_timer_second_s1_readdata                      : std_logic_vector(15 downto 0); -- timer_second:readdata -> mm_interconnect_0:timer_second_s1_readdata
	signal mm_interconnect_0_timer_second_s1_address                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_second_s1_address -> timer_second:address
	signal mm_interconnect_0_timer_second_s1_write                         : std_logic;                     -- mm_interconnect_0:timer_second_s1_write -> mm_interconnect_0_timer_second_s1_write:in
	signal mm_interconnect_0_timer_second_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_second_s1_writedata -> timer_second:writedata
	signal mm_interconnect_0_led_alarm_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:led_alarm_s1_chipselect -> led_alarm:chipselect
	signal mm_interconnect_0_led_alarm_s1_readdata                         : std_logic_vector(31 downto 0); -- led_alarm:readdata -> mm_interconnect_0:led_alarm_s1_readdata
	signal mm_interconnect_0_led_alarm_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_alarm_s1_address -> led_alarm:address
	signal mm_interconnect_0_led_alarm_s1_write                            : std_logic;                     -- mm_interconnect_0:led_alarm_s1_write -> mm_interconnect_0_led_alarm_s1_write:in
	signal mm_interconnect_0_led_alarm_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_alarm_s1_writedata -> led_alarm:writedata
	signal mm_interconnect_0_led_status_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:led_status_s1_chipselect -> led_status:chipselect
	signal mm_interconnect_0_led_status_s1_readdata                        : std_logic_vector(31 downto 0); -- led_status:readdata -> mm_interconnect_0:led_status_s1_readdata
	signal mm_interconnect_0_led_status_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_status_s1_address -> led_status:address
	signal mm_interconnect_0_led_status_s1_write                           : std_logic;                     -- mm_interconnect_0:led_status_s1_write -> mm_interconnect_0_led_status_s1_write:in
	signal mm_interconnect_0_led_status_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_status_s1_writedata -> led_status:writedata
	signal mm_interconnect_0_buttons_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:buttons_s1_chipselect -> buttons:chipselect
	signal mm_interconnect_0_buttons_s1_readdata                           : std_logic_vector(31 downto 0); -- buttons:readdata -> mm_interconnect_0:buttons_s1_readdata
	signal mm_interconnect_0_buttons_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:buttons_s1_address -> buttons:address
	signal mm_interconnect_0_buttons_s1_write                              : std_logic;                     -- mm_interconnect_0:buttons_s1_write -> mm_interconnect_0_buttons_s1_write:in
	signal mm_interconnect_0_buttons_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:buttons_s1_writedata -> buttons:writedata
	signal mm_interconnect_0_second1_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:second1_s1_chipselect -> second1:chipselect
	signal mm_interconnect_0_second1_s1_readdata                           : std_logic_vector(31 downto 0); -- second1:readdata -> mm_interconnect_0:second1_s1_readdata
	signal mm_interconnect_0_second1_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:second1_s1_address -> second1:address
	signal mm_interconnect_0_second1_s1_write                              : std_logic;                     -- mm_interconnect_0:second1_s1_write -> mm_interconnect_0_second1_s1_write:in
	signal mm_interconnect_0_second1_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:second1_s1_writedata -> second1:writedata
	signal mm_interconnect_0_minute1_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:minute1_s1_chipselect -> minute1:chipselect
	signal mm_interconnect_0_minute1_s1_readdata                           : std_logic_vector(31 downto 0); -- minute1:readdata -> mm_interconnect_0:minute1_s1_readdata
	signal mm_interconnect_0_minute1_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:minute1_s1_address -> minute1:address
	signal mm_interconnect_0_minute1_s1_write                              : std_logic;                     -- mm_interconnect_0:minute1_s1_write -> mm_interconnect_0_minute1_s1_write:in
	signal mm_interconnect_0_minute1_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:minute1_s1_writedata -> minute1:writedata
	signal mm_interconnect_0_hour1_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:hour1_s1_chipselect -> hour1:chipselect
	signal mm_interconnect_0_hour1_s1_readdata                             : std_logic_vector(31 downto 0); -- hour1:readdata -> mm_interconnect_0:hour1_s1_readdata
	signal mm_interconnect_0_hour1_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hour1_s1_address -> hour1:address
	signal mm_interconnect_0_hour1_s1_write                                : std_logic;                     -- mm_interconnect_0:hour1_s1_write -> mm_interconnect_0_hour1_s1_write:in
	signal mm_interconnect_0_hour1_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:hour1_s1_writedata -> hour1:writedata
	signal mm_interconnect_0_timer_pwm_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:timer_pwm_s1_chipselect -> timer_pwm:chipselect
	signal mm_interconnect_0_timer_pwm_s1_readdata                         : std_logic_vector(15 downto 0); -- timer_pwm:readdata -> mm_interconnect_0:timer_pwm_s1_readdata
	signal mm_interconnect_0_timer_pwm_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_pwm_s1_address -> timer_pwm:address
	signal mm_interconnect_0_timer_pwm_s1_write                            : std_logic;                     -- mm_interconnect_0:timer_pwm_s1_write -> mm_interconnect_0_timer_pwm_s1_write:in
	signal mm_interconnect_0_timer_pwm_s1_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_pwm_s1_writedata -> timer_pwm:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- timer_second:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- switches:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- buttons:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                        : std_logic;                     -- timer_pwm:irq -> irq_mapper:receiver4_irq
	signal niosii_cpu_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NiosII_CPU:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:NiosII_CPU_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_controller_reset_out_reset:in]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [NiosII_CPU:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	signal niosii_cpu_debug_reset_request_reset                            : std_logic;                     -- NiosII_CPU:debug_reset_request -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_switches_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_switches_s1_write:inv -> switches:write_n
	signal mm_interconnect_0_led_piano_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_led_piano_s1_write:inv -> led_piano:write_n
	signal mm_interconnect_0_hour0_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hour0_s1_write:inv -> hour0:write_n
	signal mm_interconnect_0_minute0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_minute0_s1_write:inv -> minute0:write_n
	signal mm_interconnect_0_second0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_second0_s1_write:inv -> second0:write_n
	signal mm_interconnect_0_timer_second_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_timer_second_s1_write:inv -> timer_second:write_n
	signal mm_interconnect_0_led_alarm_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_led_alarm_s1_write:inv -> led_alarm:write_n
	signal mm_interconnect_0_led_status_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_led_status_s1_write:inv -> led_status:write_n
	signal mm_interconnect_0_buttons_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_buttons_s1_write:inv -> buttons:write_n
	signal mm_interconnect_0_second1_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_second1_s1_write:inv -> second1:write_n
	signal mm_interconnect_0_minute1_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_minute1_s1_write:inv -> minute1:write_n
	signal mm_interconnect_0_hour1_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_hour1_s1_write:inv -> hour1:write_n
	signal mm_interconnect_0_timer_pwm_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_timer_pwm_s1_write:inv -> timer_pwm:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> NiosII_CPU:reset_n
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [buttons:reset_n, hour0:reset_n, hour1:reset_n, jtag_uart_0:rst_n, led_alarm:reset_n, led_piano:reset_n, led_status:reset_n, minute0:reset_n, minute1:reset_n, pwm:resetn, second0:reset_n, second1:reset_n, switches:reset_n, sysid_qsys_0:reset_n, timer_pwm:reset_n, timer_second:reset_n]

begin

	niosii_cpu : component qsys_system_NiosII_CPU
		port map (
			clk                                 => clk_clk,                                                  --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                 --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                       --                          .reset_req
			d_address                           => niosii_cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => niosii_cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => niosii_cpu_data_master_read,                              --                          .read
			d_readdata                          => niosii_cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => niosii_cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => niosii_cpu_data_master_write,                             --                          .write
			d_writedata                         => niosii_cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => niosii_cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => niosii_cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => niosii_cpu_instruction_master_read,                       --                          .read
			i_readdata                          => niosii_cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => niosii_cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => niosii_cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => niosii_cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => niosii_cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_niosii_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_niosii_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_niosii_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
		);

	buttons : component qsys_system_buttons
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_buttons_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_buttons_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_buttons_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_buttons_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_buttons_s1_readdata,        --                    .readdata
			in_port    => buttons_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver3_irq                      --                 irq.irq
		);

	hour0 : component qsys_system_hour0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hour0_s1_address,           --                  s1.address
			write_n    => mm_interconnect_0_hour0_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_0_hour0_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_0_hour0_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_0_hour0_s1_readdata,          --                    .readdata
			out_port   => hour0_external_connection_export              -- external_connection.export
		);

	hour1 : component qsys_system_hour0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_hour1_s1_address,           --                  s1.address
			write_n    => mm_interconnect_0_hour1_s1_write_ports_inv,   --                    .write_n
			writedata  => mm_interconnect_0_hour1_s1_writedata,         --                    .writedata
			chipselect => mm_interconnect_0_hour1_s1_chipselect,        --                    .chipselect
			readdata   => mm_interconnect_0_hour1_s1_readdata,          --                    .readdata
			out_port   => hour1_external_connection_export              -- external_connection.export
		);

	jtag_uart_0 : component qsys_system_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	led_alarm : component qsys_system_led_alarm
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_led_alarm_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_alarm_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_alarm_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_alarm_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_alarm_s1_readdata,        --                    .readdata
			out_port   => led_alarm_external_connection_export            -- external_connection.export
		);

	led_piano : component qsys_system_led_piano
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_led_piano_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_piano_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_piano_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_piano_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_piano_s1_readdata,        --                    .readdata
			out_port   => led_piano_external_connection_export            -- external_connection.export
		);

	led_status : component qsys_system_led_status
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_led_status_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_status_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_status_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_status_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_status_s1_readdata,        --                    .readdata
			out_port   => led_status_external_connection_export            -- external_connection.export
		);

	minute0 : component qsys_system_hour0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_minute0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_minute0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_minute0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_minute0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_minute0_s1_readdata,        --                    .readdata
			out_port   => minute0_external_connection_export            -- external_connection.export
		);

	minute1 : component qsys_system_hour0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_minute1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_minute1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_minute1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_minute1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_minute1_s1_readdata,        --                    .readdata
			out_port   => minute1_external_connection_export            -- external_connection.export
		);

	onchip_memory : component qsys_system_onchip_memory
		port map (
			clk        => clk_clk,                                       --   clk1.clk
			address    => mm_interconnect_0_onchip_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                            -- (terminated)
		);

	pwm : component pwm_avalon_interface
		generic map (
			clock_divide_reg_init => "0000000000000000000000000000000000",
			duty_cycle_reg_init   => "0000000000000000000000000000000000"
		)
		port map (
			clk                => clk_clk,                                        --         clock.clk
			pwm_out            => pwm_external_connection_export,                 --       pwm_out.export
			resetn             => rst_controller_001_reset_out_reset_ports_inv,   --        resetn.reset_n
			avalon_chip_select => mm_interconnect_0_pwm_control_slave_chipselect, -- control_slave.chipselect
			address            => mm_interconnect_0_pwm_control_slave_address,    --              .address
			write              => mm_interconnect_0_pwm_control_slave_write,      --              .write
			write_data         => mm_interconnect_0_pwm_control_slave_writedata,  --              .writedata
			read               => mm_interconnect_0_pwm_control_slave_read,       --              .read
			read_data          => mm_interconnect_0_pwm_control_slave_readdata    --              .readdata
		);

	second0 : component qsys_system_hour0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_second0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_second0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_second0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_second0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_second0_s1_readdata,        --                    .readdata
			out_port   => second0_external_connection_export            -- external_connection.export
		);

	second1 : component qsys_system_hour0
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_second1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_second1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_second1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_second1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_second1_s1_readdata,        --                    .readdata
			out_port   => second1_external_connection_export            -- external_connection.export
		);

	switches : component qsys_system_switches
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_switches_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_switches_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_switches_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_switches_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_switches_s1_readdata,        --                    .readdata
			in_port    => switches_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                       --                 irq.irq
		);

	sysid_qsys_0 : component qsys_system_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,            --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_pwm : component qsys_system_timer_pwm
		port map (
			clk        => clk_clk,                                        --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_pwm_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_pwm_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_pwm_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_pwm_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_pwm_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver4_irq                        --   irq.irq
		);

	timer_second : component qsys_system_timer_second
		port map (
			clk        => clk_clk,                                           --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,      -- reset.reset_n
			address    => mm_interconnect_0_timer_second_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_second_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_second_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_second_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_second_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                           --   irq.irq
		);

	mm_interconnect_0 : component qsys_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                 => clk_clk,                                                     --                               clk_0_clk.clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                          -- jtag_uart_0_reset_reset_bridge_in_reset.reset
			NiosII_CPU_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                              --  NiosII_CPU_reset_reset_bridge_in_reset.reset
			NiosII_CPU_data_master_address                => niosii_cpu_data_master_address,                              --                  NiosII_CPU_data_master.address
			NiosII_CPU_data_master_waitrequest            => niosii_cpu_data_master_waitrequest,                          --                                        .waitrequest
			NiosII_CPU_data_master_byteenable             => niosii_cpu_data_master_byteenable,                           --                                        .byteenable
			NiosII_CPU_data_master_read                   => niosii_cpu_data_master_read,                                 --                                        .read
			NiosII_CPU_data_master_readdata               => niosii_cpu_data_master_readdata,                             --                                        .readdata
			NiosII_CPU_data_master_write                  => niosii_cpu_data_master_write,                                --                                        .write
			NiosII_CPU_data_master_writedata              => niosii_cpu_data_master_writedata,                            --                                        .writedata
			NiosII_CPU_data_master_debugaccess            => niosii_cpu_data_master_debugaccess,                          --                                        .debugaccess
			NiosII_CPU_instruction_master_address         => niosii_cpu_instruction_master_address,                       --           NiosII_CPU_instruction_master.address
			NiosII_CPU_instruction_master_waitrequest     => niosii_cpu_instruction_master_waitrequest,                   --                                        .waitrequest
			NiosII_CPU_instruction_master_read            => niosii_cpu_instruction_master_read,                          --                                        .read
			NiosII_CPU_instruction_master_readdata        => niosii_cpu_instruction_master_readdata,                      --                                        .readdata
			NiosII_CPU_instruction_master_readdatavalid   => niosii_cpu_instruction_master_readdatavalid,                 --                                        .readdatavalid
			buttons_s1_address                            => mm_interconnect_0_buttons_s1_address,                        --                              buttons_s1.address
			buttons_s1_write                              => mm_interconnect_0_buttons_s1_write,                          --                                        .write
			buttons_s1_readdata                           => mm_interconnect_0_buttons_s1_readdata,                       --                                        .readdata
			buttons_s1_writedata                          => mm_interconnect_0_buttons_s1_writedata,                      --                                        .writedata
			buttons_s1_chipselect                         => mm_interconnect_0_buttons_s1_chipselect,                     --                                        .chipselect
			hour0_s1_address                              => mm_interconnect_0_hour0_s1_address,                          --                                hour0_s1.address
			hour0_s1_write                                => mm_interconnect_0_hour0_s1_write,                            --                                        .write
			hour0_s1_readdata                             => mm_interconnect_0_hour0_s1_readdata,                         --                                        .readdata
			hour0_s1_writedata                            => mm_interconnect_0_hour0_s1_writedata,                        --                                        .writedata
			hour0_s1_chipselect                           => mm_interconnect_0_hour0_s1_chipselect,                       --                                        .chipselect
			hour1_s1_address                              => mm_interconnect_0_hour1_s1_address,                          --                                hour1_s1.address
			hour1_s1_write                                => mm_interconnect_0_hour1_s1_write,                            --                                        .write
			hour1_s1_readdata                             => mm_interconnect_0_hour1_s1_readdata,                         --                                        .readdata
			hour1_s1_writedata                            => mm_interconnect_0_hour1_s1_writedata,                        --                                        .writedata
			hour1_s1_chipselect                           => mm_interconnect_0_hour1_s1_chipselect,                       --                                        .chipselect
			jtag_uart_0_avalon_jtag_slave_address         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --           jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                        .write
			jtag_uart_0_avalon_jtag_slave_read            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                        .read
			jtag_uart_0_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                        .readdata
			jtag_uart_0_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                        .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                        .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                        .chipselect
			led_alarm_s1_address                          => mm_interconnect_0_led_alarm_s1_address,                      --                            led_alarm_s1.address
			led_alarm_s1_write                            => mm_interconnect_0_led_alarm_s1_write,                        --                                        .write
			led_alarm_s1_readdata                         => mm_interconnect_0_led_alarm_s1_readdata,                     --                                        .readdata
			led_alarm_s1_writedata                        => mm_interconnect_0_led_alarm_s1_writedata,                    --                                        .writedata
			led_alarm_s1_chipselect                       => mm_interconnect_0_led_alarm_s1_chipselect,                   --                                        .chipselect
			led_piano_s1_address                          => mm_interconnect_0_led_piano_s1_address,                      --                            led_piano_s1.address
			led_piano_s1_write                            => mm_interconnect_0_led_piano_s1_write,                        --                                        .write
			led_piano_s1_readdata                         => mm_interconnect_0_led_piano_s1_readdata,                     --                                        .readdata
			led_piano_s1_writedata                        => mm_interconnect_0_led_piano_s1_writedata,                    --                                        .writedata
			led_piano_s1_chipselect                       => mm_interconnect_0_led_piano_s1_chipselect,                   --                                        .chipselect
			led_status_s1_address                         => mm_interconnect_0_led_status_s1_address,                     --                           led_status_s1.address
			led_status_s1_write                           => mm_interconnect_0_led_status_s1_write,                       --                                        .write
			led_status_s1_readdata                        => mm_interconnect_0_led_status_s1_readdata,                    --                                        .readdata
			led_status_s1_writedata                       => mm_interconnect_0_led_status_s1_writedata,                   --                                        .writedata
			led_status_s1_chipselect                      => mm_interconnect_0_led_status_s1_chipselect,                  --                                        .chipselect
			minute0_s1_address                            => mm_interconnect_0_minute0_s1_address,                        --                              minute0_s1.address
			minute0_s1_write                              => mm_interconnect_0_minute0_s1_write,                          --                                        .write
			minute0_s1_readdata                           => mm_interconnect_0_minute0_s1_readdata,                       --                                        .readdata
			minute0_s1_writedata                          => mm_interconnect_0_minute0_s1_writedata,                      --                                        .writedata
			minute0_s1_chipselect                         => mm_interconnect_0_minute0_s1_chipselect,                     --                                        .chipselect
			minute1_s1_address                            => mm_interconnect_0_minute1_s1_address,                        --                              minute1_s1.address
			minute1_s1_write                              => mm_interconnect_0_minute1_s1_write,                          --                                        .write
			minute1_s1_readdata                           => mm_interconnect_0_minute1_s1_readdata,                       --                                        .readdata
			minute1_s1_writedata                          => mm_interconnect_0_minute1_s1_writedata,                      --                                        .writedata
			minute1_s1_chipselect                         => mm_interconnect_0_minute1_s1_chipselect,                     --                                        .chipselect
			NiosII_CPU_debug_mem_slave_address            => mm_interconnect_0_niosii_cpu_debug_mem_slave_address,        --              NiosII_CPU_debug_mem_slave.address
			NiosII_CPU_debug_mem_slave_write              => mm_interconnect_0_niosii_cpu_debug_mem_slave_write,          --                                        .write
			NiosII_CPU_debug_mem_slave_read               => mm_interconnect_0_niosii_cpu_debug_mem_slave_read,           --                                        .read
			NiosII_CPU_debug_mem_slave_readdata           => mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata,       --                                        .readdata
			NiosII_CPU_debug_mem_slave_writedata          => mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata,      --                                        .writedata
			NiosII_CPU_debug_mem_slave_byteenable         => mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable,     --                                        .byteenable
			NiosII_CPU_debug_mem_slave_waitrequest        => mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest,    --                                        .waitrequest
			NiosII_CPU_debug_mem_slave_debugaccess        => mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess,    --                                        .debugaccess
			onchip_memory_s1_address                      => mm_interconnect_0_onchip_memory_s1_address,                  --                        onchip_memory_s1.address
			onchip_memory_s1_write                        => mm_interconnect_0_onchip_memory_s1_write,                    --                                        .write
			onchip_memory_s1_readdata                     => mm_interconnect_0_onchip_memory_s1_readdata,                 --                                        .readdata
			onchip_memory_s1_writedata                    => mm_interconnect_0_onchip_memory_s1_writedata,                --                                        .writedata
			onchip_memory_s1_byteenable                   => mm_interconnect_0_onchip_memory_s1_byteenable,               --                                        .byteenable
			onchip_memory_s1_chipselect                   => mm_interconnect_0_onchip_memory_s1_chipselect,               --                                        .chipselect
			onchip_memory_s1_clken                        => mm_interconnect_0_onchip_memory_s1_clken,                    --                                        .clken
			pwm_control_slave_address                     => mm_interconnect_0_pwm_control_slave_address,                 --                       pwm_control_slave.address
			pwm_control_slave_write                       => mm_interconnect_0_pwm_control_slave_write,                   --                                        .write
			pwm_control_slave_read                        => mm_interconnect_0_pwm_control_slave_read,                    --                                        .read
			pwm_control_slave_readdata                    => mm_interconnect_0_pwm_control_slave_readdata,                --                                        .readdata
			pwm_control_slave_writedata                   => mm_interconnect_0_pwm_control_slave_writedata,               --                                        .writedata
			pwm_control_slave_chipselect                  => mm_interconnect_0_pwm_control_slave_chipselect,              --                                        .chipselect
			second0_s1_address                            => mm_interconnect_0_second0_s1_address,                        --                              second0_s1.address
			second0_s1_write                              => mm_interconnect_0_second0_s1_write,                          --                                        .write
			second0_s1_readdata                           => mm_interconnect_0_second0_s1_readdata,                       --                                        .readdata
			second0_s1_writedata                          => mm_interconnect_0_second0_s1_writedata,                      --                                        .writedata
			second0_s1_chipselect                         => mm_interconnect_0_second0_s1_chipselect,                     --                                        .chipselect
			second1_s1_address                            => mm_interconnect_0_second1_s1_address,                        --                              second1_s1.address
			second1_s1_write                              => mm_interconnect_0_second1_s1_write,                          --                                        .write
			second1_s1_readdata                           => mm_interconnect_0_second1_s1_readdata,                       --                                        .readdata
			second1_s1_writedata                          => mm_interconnect_0_second1_s1_writedata,                      --                                        .writedata
			second1_s1_chipselect                         => mm_interconnect_0_second1_s1_chipselect,                     --                                        .chipselect
			switches_s1_address                           => mm_interconnect_0_switches_s1_address,                       --                             switches_s1.address
			switches_s1_write                             => mm_interconnect_0_switches_s1_write,                         --                                        .write
			switches_s1_readdata                          => mm_interconnect_0_switches_s1_readdata,                      --                                        .readdata
			switches_s1_writedata                         => mm_interconnect_0_switches_s1_writedata,                     --                                        .writedata
			switches_s1_chipselect                        => mm_interconnect_0_switches_s1_chipselect,                    --                                        .chipselect
			sysid_qsys_0_control_slave_address            => mm_interconnect_0_sysid_qsys_0_control_slave_address,        --              sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata           => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,       --                                        .readdata
			timer_pwm_s1_address                          => mm_interconnect_0_timer_pwm_s1_address,                      --                            timer_pwm_s1.address
			timer_pwm_s1_write                            => mm_interconnect_0_timer_pwm_s1_write,                        --                                        .write
			timer_pwm_s1_readdata                         => mm_interconnect_0_timer_pwm_s1_readdata,                     --                                        .readdata
			timer_pwm_s1_writedata                        => mm_interconnect_0_timer_pwm_s1_writedata,                    --                                        .writedata
			timer_pwm_s1_chipselect                       => mm_interconnect_0_timer_pwm_s1_chipselect,                   --                                        .chipselect
			timer_second_s1_address                       => mm_interconnect_0_timer_second_s1_address,                   --                         timer_second_s1.address
			timer_second_s1_write                         => mm_interconnect_0_timer_second_s1_write,                     --                                        .write
			timer_second_s1_readdata                      => mm_interconnect_0_timer_second_s1_readdata,                  --                                        .readdata
			timer_second_s1_writedata                     => mm_interconnect_0_timer_second_s1_writedata,                 --                                        .writedata
			timer_second_s1_chipselect                    => mm_interconnect_0_timer_second_s1_chipselect                 --                                        .chipselect
		);

	irq_mapper : component qsys_system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			sender_irq    => niosii_cpu_irq_irq              --    sender.irq
		);

	rst_controller : component qsys_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,              -- reset_in0.reset
			reset_in1      => niosii_cpu_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                              --       clk.clk
			reset_out      => rst_controller_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_001 : component qsys_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_switches_s1_write_ports_inv <= not mm_interconnect_0_switches_s1_write;

	mm_interconnect_0_led_piano_s1_write_ports_inv <= not mm_interconnect_0_led_piano_s1_write;

	mm_interconnect_0_hour0_s1_write_ports_inv <= not mm_interconnect_0_hour0_s1_write;

	mm_interconnect_0_minute0_s1_write_ports_inv <= not mm_interconnect_0_minute0_s1_write;

	mm_interconnect_0_second0_s1_write_ports_inv <= not mm_interconnect_0_second0_s1_write;

	mm_interconnect_0_timer_second_s1_write_ports_inv <= not mm_interconnect_0_timer_second_s1_write;

	mm_interconnect_0_led_alarm_s1_write_ports_inv <= not mm_interconnect_0_led_alarm_s1_write;

	mm_interconnect_0_led_status_s1_write_ports_inv <= not mm_interconnect_0_led_status_s1_write;

	mm_interconnect_0_buttons_s1_write_ports_inv <= not mm_interconnect_0_buttons_s1_write;

	mm_interconnect_0_second1_s1_write_ports_inv <= not mm_interconnect_0_second1_s1_write;

	mm_interconnect_0_minute1_s1_write_ports_inv <= not mm_interconnect_0_minute1_s1_write;

	mm_interconnect_0_hour1_s1_write_ports_inv <= not mm_interconnect_0_hour1_s1_write;

	mm_interconnect_0_timer_pwm_s1_write_ports_inv <= not mm_interconnect_0_timer_pwm_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of qsys_system
